LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY distance2clkdivisor IS
   PORT(
			clk            :  IN    STD_LOGIC;                                
			reset          :  IN    STD_LOGIC; 
			distance       :  IN    STD_LOGIC_VECTOR(12 DOWNTO 0);                           
			divisor        :  OUT   natural
		  );  
END distance2clkdivisor;

ARCHITECTURE behavior OF distance2clkdivisor IS

type array_1d is array (0 to 4095) of integer;

constant d2d_LUT : array_1d := ( 
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	3	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	4	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	5	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	6	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	7	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	8	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	9	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	10	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	15	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	20	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	30	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	50	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	100	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	),
(	200	)
);

begin

divisor <= d2d_LUT(to_integer(unsigned(distance)));
							
end behavior;
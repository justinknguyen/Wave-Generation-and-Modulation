LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY distance2cycle IS
   PORT(
			clk            :  IN    STD_LOGIC;                                
			reset          :  IN    STD_LOGIC; 
			distance       :  IN    STD_LOGIC_VECTOR(12 DOWNTO 0);                           
			cycle	         :  OUT   STD_LOGIC_VECTOR(12 DOWNTO 0)
		  );  
END distance2cycle;

ARCHITECTURE behavior OF distance2cycle IS

type array_1d is array (0 to 4095) of integer;

constant d2c_LUT : array_1d := ( 
(	8190	),
(	8180	),
(	8180	),
(	8180	),
(	8170	),
(	8170	),
(	8170	),
(	8170	),
(	8160	),
(	8160	),
(	8160	),
(	8150	),
(	8150	),
(	8150	),
(	8140	),
(	8140	),
(	8140	),
(	8140	),
(	8130	),
(	8130	),
(	8130	),
(	8120	),
(	8120	),
(	8120	),
(	8120	),
(	8110	),
(	8110	),
(	8110	),
(	8100	),
(	8100	),
(	8100	),
(	8090	),
(	8090	),
(	8090	),
(	8090	),
(	8080	),
(	8080	),
(	8080	),
(	8070	),
(	8070	),
(	8070	),
(	8070	),
(	8060	),
(	8060	),
(	8060	),
(	8050	),
(	8050	),
(	8050	),
(	8040	),
(	8040	),
(	8040	),
(	8040	),
(	8030	),
(	8030	),
(	8030	),
(	8020	),
(	8020	),
(	8020	),
(	8020	),
(	8010	),
(	8010	),
(	8010	),
(	8000	),
(	8000	),
(	8000	),
(	7990	),
(	7990	),
(	7990	),
(	7990	),
(	7980	),
(	7980	),
(	7980	),
(	7970	),
(	7970	),
(	7970	),
(	7970	),
(	7960	),
(	7960	),
(	7960	),
(	7950	),
(	7950	),
(	7950	),
(	7940	),
(	7940	),
(	7940	),
(	7940	),
(	7930	),
(	7930	),
(	7930	),
(	7920	),
(	7920	),
(	7920	),
(	7920	),
(	7910	),
(	7910	),
(	7910	),
(	7900	),
(	7900	),
(	7900	),
(	7890	),
(	7890	),
(	7890	),
(	7890	),
(	7880	),
(	7880	),
(	7880	),
(	7870	),
(	7870	),
(	7870	),
(	7870	),
(	7860	),
(	7860	),
(	7860	),
(	7850	),
(	7850	),
(	7850	),
(	7840	),
(	7840	),
(	7840	),
(	7840	),
(	7830	),
(	7830	),
(	7830	),
(	7820	),
(	7820	),
(	7820	),
(	7820	),
(	7810	),
(	7810	),
(	7810	),
(	7800	),
(	7800	),
(	7800	),
(	7790	),
(	7790	),
(	7790	),
(	7790	),
(	7780	),
(	7780	),
(	7780	),
(	7770	),
(	7770	),
(	7770	),
(	7770	),
(	7760	),
(	7760	),
(	7760	),
(	7750	),
(	7750	),
(	7750	),
(	7750	),
(	7740	),
(	7740	),
(	7740	),
(	7730	),
(	7730	),
(	7730	),
(	7720	),
(	7720	),
(	7720	),
(	7720	),
(	7710	),
(	7710	),
(	7710	),
(	7700	),
(	7700	),
(	7700	),
(	7700	),
(	7690	),
(	7690	),
(	7690	),
(	7680	),
(	7680	),
(	7680	),
(	7670	),
(	7670	),
(	7670	),
(	7670	),
(	7660	),
(	7660	),
(	7660	),
(	7650	),
(	7650	),
(	7650	),
(	7650	),
(	7640	),
(	7640	),
(	7640	),
(	7630	),
(	7630	),
(	7630	),
(	7620	),
(	7620	),
(	7620	),
(	7620	),
(	7610	),
(	7610	),
(	7610	),
(	7600	),
(	7600	),
(	7600	),
(	7600	),
(	7590	),
(	7590	),
(	7590	),
(	7580	),
(	7580	),
(	7580	),
(	7570	),
(	7570	),
(	7570	),
(	7570	),
(	7560	),
(	7560	),
(	7560	),
(	7550	),
(	7550	),
(	7550	),
(	7550	),
(	7540	),
(	7540	),
(	7540	),
(	7530	),
(	7530	),
(	7530	),
(	7520	),
(	7520	),
(	7520	),
(	7520	),
(	7510	),
(	7510	),
(	7510	),
(	7500	),
(	7500	),
(	7500	),
(	7500	),
(	7490	),
(	7490	),
(	7490	),
(	7480	),
(	7480	),
(	7480	),
(	7470	),
(	7470	),
(	7470	),
(	7470	),
(	7460	),
(	7460	),
(	7460	),
(	7450	),
(	7450	),
(	7450	),
(	7450	),
(	7440	),
(	7440	),
(	7440	),
(	7430	),
(	7430	),
(	7430	),
(	7420	),
(	7420	),
(	7420	),
(	7420	),
(	7410	),
(	7410	),
(	7410	),
(	7400	),
(	7400	),
(	7400	),
(	7400	),
(	7390	),
(	7390	),
(	7390	),
(	7380	),
(	7380	),
(	7380	),
(	7370	),
(	7370	),
(	7370	),
(	7370	),
(	7360	),
(	7360	),
(	7360	),
(	7350	),
(	7350	),
(	7350	),
(	7350	),
(	7340	),
(	7340	),
(	7340	),
(	7330	),
(	7330	),
(	7330	),
(	7320	),
(	7320	),
(	7320	),
(	7320	),
(	7310	),
(	7310	),
(	7310	),
(	7300	),
(	7300	),
(	7300	),
(	7300	),
(	7290	),
(	7290	),
(	7290	),
(	7280	),
(	7280	),
(	7280	),
(	7270	),
(	7270	),
(	7270	),
(	7270	),
(	7260	),
(	7260	),
(	7260	),
(	7250	),
(	7250	),
(	7250	),
(	7250	),
(	7240	),
(	7240	),
(	7240	),
(	7230	),
(	7230	),
(	7230	),
(	7220	),
(	7220	),
(	7220	),
(	7220	),
(	7210	),
(	7210	),
(	7210	),
(	7200	),
(	7200	),
(	7200	),
(	7200	),
(	7190	),
(	7190	),
(	7190	),
(	7180	),
(	7180	),
(	7180	),
(	7170	),
(	7170	),
(	7170	),
(	7170	),
(	7160	),
(	7160	),
(	7160	),
(	7150	),
(	7150	),
(	7150	),
(	7150	),
(	7140	),
(	7140	),
(	7140	),
(	7130	),
(	7130	),
(	7130	),
(	7120	),
(	7120	),
(	7120	),
(	7120	),
(	7110	),
(	7110	),
(	7110	),
(	7100	),
(	7100	),
(	7100	),
(	7100	),
(	7090	),
(	7090	),
(	7090	),
(	7080	),
(	7080	),
(	7080	),
(	7070	),
(	7070	),
(	7070	),
(	7070	),
(	7060	),
(	7060	),
(	7060	),
(	7050	),
(	7050	),
(	7050	),
(	7050	),
(	7040	),
(	7040	),
(	7040	),
(	7030	),
(	7030	),
(	7030	),
(	7020	),
(	7020	),
(	7020	),
(	7020	),
(	7010	),
(	7010	),
(	7010	),
(	7000	),
(	7000	),
(	7000	),
(	7000	),
(	6990	),
(	6990	),
(	6990	),
(	6980	),
(	6980	),
(	6980	),
(	6970	),
(	6970	),
(	6970	),
(	6970	),
(	6960	),
(	6960	),
(	6960	),
(	6950	),
(	6950	),
(	6950	),
(	6950	),
(	6940	),
(	6940	),
(	6940	),
(	6930	),
(	6930	),
(	6930	),
(	6920	),
(	6920	),
(	6920	),
(	6920	),
(	6910	),
(	6910	),
(	6910	),
(	6900	),
(	6900	),
(	6900	),
(	6900	),
(	6890	),
(	6890	),
(	6890	),
(	6880	),
(	6880	),
(	6880	),
(	6870	),
(	6870	),
(	6870	),
(	6870	),
(	6860	),
(	6860	),
(	6860	),
(	6850	),
(	6850	),
(	6850	),
(	6850	),
(	6840	),
(	6840	),
(	6840	),
(	6830	),
(	6830	),
(	6830	),
(	6820	),
(	6820	),
(	6820	),
(	6820	),
(	6810	),
(	6810	),
(	6810	),
(	6800	),
(	6800	),
(	6800	),
(	6800	),
(	6790	),
(	6790	),
(	6790	),
(	6780	),
(	6780	),
(	6780	),
(	6770	),
(	6770	),
(	6770	),
(	6770	),
(	6760	),
(	6760	),
(	6760	),
(	6750	),
(	6750	),
(	6750	),
(	6750	),
(	6740	),
(	6740	),
(	6740	),
(	6730	),
(	6730	),
(	6730	),
(	6720	),
(	6720	),
(	6720	),
(	6720	),
(	6710	),
(	6710	),
(	6710	),
(	6700	),
(	6700	),
(	6700	),
(	6700	),
(	6690	),
(	6690	),
(	6690	),
(	6680	),
(	6680	),
(	6680	),
(	6670	),
(	6670	),
(	6670	),
(	6670	),
(	6660	),
(	6660	),
(	6660	),
(	6650	),
(	6650	),
(	6650	),
(	6650	),
(	6640	),
(	6640	),
(	6640	),
(	6630	),
(	6630	),
(	6630	),
(	6620	),
(	6620	),
(	6620	),
(	6620	),
(	6610	),
(	6610	),
(	6610	),
(	6600	),
(	6600	),
(	6600	),
(	6600	),
(	6590	),
(	6590	),
(	6590	),
(	6580	),
(	6580	),
(	6580	),
(	6570	),
(	6570	),
(	6570	),
(	6570	),
(	6560	),
(	6560	),
(	6560	),
(	6550	),
(	6550	),
(	6550	),
(	6550	),
(	6540	),
(	6540	),
(	6540	),
(	6530	),
(	6530	),
(	6530	),
(	6520	),
(	6520	),
(	6520	),
(	6520	),
(	6510	),
(	6510	),
(	6510	),
(	6500	),
(	6500	),
(	6500	),
(	6500	),
(	6490	),
(	6490	),
(	6490	),
(	6480	),
(	6480	),
(	6480	),
(	6470	),
(	6470	),
(	6470	),
(	6470	),
(	6460	),
(	6460	),
(	6460	),
(	6450	),
(	6450	),
(	6450	),
(	6450	),
(	6440	),
(	6440	),
(	6440	),
(	6430	),
(	6430	),
(	6430	),
(	6420	),
(	6420	),
(	6420	),
(	6420	),
(	6410	),
(	6410	),
(	6410	),
(	6400	),
(	6400	),
(	6400	),
(	6400	),
(	6390	),
(	6390	),
(	6390	),
(	6380	),
(	6380	),
(	6380	),
(	6380	),
(	6370	),
(	6370	),
(	6370	),
(	6360	),
(	6360	),
(	6360	),
(	6350	),
(	6350	),
(	6350	),
(	6350	),
(	6340	),
(	6340	),
(	6340	),
(	6330	),
(	6330	),
(	6330	),
(	6330	),
(	6320	),
(	6320	),
(	6320	),
(	6310	),
(	6310	),
(	6310	),
(	6300	),
(	6300	),
(	6300	),
(	6300	),
(	6290	),
(	6290	),
(	6290	),
(	6280	),
(	6280	),
(	6280	),
(	6280	),
(	6270	),
(	6270	),
(	6270	),
(	6260	),
(	6260	),
(	6260	),
(	6250	),
(	6250	),
(	6250	),
(	6250	),
(	6240	),
(	6240	),
(	6240	),
(	6230	),
(	6230	),
(	6230	),
(	6230	),
(	6220	),
(	6220	),
(	6220	),
(	6210	),
(	6210	),
(	6210	),
(	6200	),
(	6200	),
(	6200	),
(	6200	),
(	6190	),
(	6190	),
(	6190	),
(	6180	),
(	6180	),
(	6180	),
(	6180	),
(	6170	),
(	6170	),
(	6170	),
(	6160	),
(	6160	),
(	6160	),
(	6150	),
(	6150	),
(	6150	),
(	6150	),
(	6140	),
(	6140	),
(	6140	),
(	6130	),
(	6130	),
(	6130	),
(	6130	),
(	6120	),
(	6120	),
(	6120	),
(	6110	),
(	6110	),
(	6110	),
(	6100	),
(	6100	),
(	6100	),
(	6100	),
(	6090	),
(	6090	),
(	6090	),
(	6080	),
(	6080	),
(	6080	),
(	6080	),
(	6070	),
(	6070	),
(	6070	),
(	6060	),
(	6060	),
(	6060	),
(	6050	),
(	6050	),
(	6050	),
(	6050	),
(	6040	),
(	6040	),
(	6040	),
(	6030	),
(	6030	),
(	6030	),
(	6030	),
(	6020	),
(	6020	),
(	6020	),
(	6010	),
(	6010	),
(	6010	),
(	6000	),
(	6000	),
(	6000	),
(	6000	),
(	5990	),
(	5990	),
(	5990	),
(	5980	),
(	5980	),
(	5980	),
(	5980	),
(	5970	),
(	5970	),
(	5970	),
(	5960	),
(	5960	),
(	5960	),
(	5950	),
(	5950	),
(	5950	),
(	5950	),
(	5940	),
(	5940	),
(	5940	),
(	5930	),
(	5930	),
(	5930	),
(	5930	),
(	5920	),
(	5920	),
(	5920	),
(	5910	),
(	5910	),
(	5910	),
(	5900	),
(	5900	),
(	5900	),
(	5900	),
(	5890	),
(	5890	),
(	5890	),
(	5880	),
(	5880	),
(	5880	),
(	5880	),
(	5870	),
(	5870	),
(	5870	),
(	5860	),
(	5860	),
(	5860	),
(	5850	),
(	5850	),
(	5850	),
(	5850	),
(	5840	),
(	5840	),
(	5840	),
(	5830	),
(	5830	),
(	5830	),
(	5830	),
(	5820	),
(	5820	),
(	5820	),
(	5810	),
(	5810	),
(	5810	),
(	5800	),
(	5800	),
(	5800	),
(	5800	),
(	5790	),
(	5790	),
(	5790	),
(	5780	),
(	5780	),
(	5780	),
(	5780	),
(	5770	),
(	5770	),
(	5770	),
(	5760	),
(	5760	),
(	5760	),
(	5750	),
(	5750	),
(	5750	),
(	5750	),
(	5740	),
(	5740	),
(	5740	),
(	5730	),
(	5730	),
(	5730	),
(	5730	),
(	5720	),
(	5720	),
(	5720	),
(	5710	),
(	5710	),
(	5710	),
(	5700	),
(	5700	),
(	5700	),
(	5700	),
(	5690	),
(	5690	),
(	5690	),
(	5680	),
(	5680	),
(	5680	),
(	5680	),
(	5670	),
(	5670	),
(	5670	),
(	5660	),
(	5660	),
(	5660	),
(	5650	),
(	5650	),
(	5650	),
(	5650	),
(	5640	),
(	5640	),
(	5640	),
(	5630	),
(	5630	),
(	5630	),
(	5630	),
(	5620	),
(	5620	),
(	5620	),
(	5610	),
(	5610	),
(	5610	),
(	5600	),
(	5600	),
(	5600	),
(	5600	),
(	5590	),
(	5590	),
(	5590	),
(	5580	),
(	5580	),
(	5580	),
(	5580	),
(	5570	),
(	5570	),
(	5570	),
(	5560	),
(	5560	),
(	5560	),
(	5550	),
(	5550	),
(	5550	),
(	5550	),
(	5540	),
(	5540	),
(	5540	),
(	5530	),
(	5530	),
(	5530	),
(	5530	),
(	5520	),
(	5520	),
(	5520	),
(	5510	),
(	5510	),
(	5510	),
(	5500	),
(	5500	),
(	5500	),
(	5500	),
(	5490	),
(	5490	),
(	5490	),
(	5480	),
(	5480	),
(	5480	),
(	5480	),
(	5470	),
(	5470	),
(	5470	),
(	5460	),
(	5460	),
(	5460	),
(	5450	),
(	5450	),
(	5450	),
(	5450	),
(	5440	),
(	5440	),
(	5440	),
(	5430	),
(	5430	),
(	5430	),
(	5430	),
(	5420	),
(	5420	),
(	5420	),
(	5410	),
(	5410	),
(	5410	),
(	5400	),
(	5400	),
(	5400	),
(	5400	),
(	5390	),
(	5390	),
(	5390	),
(	5380	),
(	5380	),
(	5380	),
(	5380	),
(	5370	),
(	5370	),
(	5370	),
(	5360	),
(	5360	),
(	5360	),
(	5350	),
(	5350	),
(	5350	),
(	5350	),
(	5340	),
(	5340	),
(	5340	),
(	5330	),
(	5330	),
(	5330	),
(	5330	),
(	5320	),
(	5320	),
(	5320	),
(	5310	),
(	5310	),
(	5310	),
(	5300	),
(	5300	),
(	5300	),
(	5300	),
(	5290	),
(	5290	),
(	5290	),
(	5280	),
(	5280	),
(	5280	),
(	5280	),
(	5270	),
(	5270	),
(	5270	),
(	5260	),
(	5260	),
(	5260	),
(	5250	),
(	5250	),
(	5250	),
(	5250	),
(	5240	),
(	5240	),
(	5240	),
(	5230	),
(	5230	),
(	5230	),
(	5230	),
(	5220	),
(	5220	),
(	5220	),
(	5210	),
(	5210	),
(	5210	),
(	5200	),
(	5200	),
(	5200	),
(	5200	),
(	5190	),
(	5190	),
(	5190	),
(	5180	),
(	5180	),
(	5180	),
(	5180	),
(	5170	),
(	5170	),
(	5170	),
(	5160	),
(	5160	),
(	5160	),
(	5150	),
(	5150	),
(	5150	),
(	5150	),
(	5140	),
(	5140	),
(	5140	),
(	5130	),
(	5130	),
(	5130	),
(	5130	),
(	5120	),
(	5120	),
(	5120	),
(	5110	),
(	5110	),
(	5110	),
(	5100	),
(	5100	),
(	5100	),
(	5100	),
(	5090	),
(	5090	),
(	5090	),
(	5080	),
(	5080	),
(	5080	),
(	5080	),
(	5070	),
(	5070	),
(	5070	),
(	5060	),
(	5060	),
(	5060	),
(	5050	),
(	5050	),
(	5050	),
(	5050	),
(	5040	),
(	5040	),
(	5040	),
(	5030	),
(	5030	),
(	5030	),
(	5030	),
(	5020	),
(	5020	),
(	5020	),
(	5010	),
(	5010	),
(	5010	),
(	5010	),
(	5000	),
(	5000	),
(	5000	),
(	4990	),
(	4990	),
(	4990	),
(	4980	),
(	4980	),
(	4980	),
(	4980	),
(	4970	),
(	4970	),
(	4970	),
(	4960	),
(	4960	),
(	4960	),
(	4960	),
(	4950	),
(	4950	),
(	4950	),
(	4940	),
(	4940	),
(	4940	),
(	4930	),
(	4930	),
(	4930	),
(	4930	),
(	4920	),
(	4920	),
(	4920	),
(	4910	),
(	4910	),
(	4910	),
(	4910	),
(	4900	),
(	4900	),
(	4900	),
(	4890	),
(	4890	),
(	4890	),
(	4880	),
(	4880	),
(	4880	),
(	4880	),
(	4870	),
(	4870	),
(	4870	),
(	4860	),
(	4860	),
(	4860	),
(	4860	),
(	4850	),
(	4850	),
(	4850	),
(	4840	),
(	4840	),
(	4840	),
(	4830	),
(	4830	),
(	4830	),
(	4830	),
(	4820	),
(	4820	),
(	4820	),
(	4810	),
(	4810	),
(	4810	),
(	4810	),
(	4800	),
(	4800	),
(	4800	),
(	4790	),
(	4790	),
(	4790	),
(	4780	),
(	4780	),
(	4780	),
(	4780	),
(	4770	),
(	4770	),
(	4770	),
(	4760	),
(	4760	),
(	4760	),
(	4760	),
(	4750	),
(	4750	),
(	4750	),
(	4740	),
(	4740	),
(	4740	),
(	4730	),
(	4730	),
(	4730	),
(	4730	),
(	4720	),
(	4720	),
(	4720	),
(	4710	),
(	4710	),
(	4710	),
(	4710	),
(	4700	),
(	4700	),
(	4700	),
(	4690	),
(	4690	),
(	4690	),
(	4680	),
(	4680	),
(	4680	),
(	4680	),
(	4670	),
(	4670	),
(	4670	),
(	4660	),
(	4660	),
(	4660	),
(	4660	),
(	4650	),
(	4650	),
(	4650	),
(	4640	),
(	4640	),
(	4640	),
(	4630	),
(	4630	),
(	4630	),
(	4630	),
(	4620	),
(	4620	),
(	4620	),
(	4610	),
(	4610	),
(	4610	),
(	4610	),
(	4600	),
(	4600	),
(	4600	),
(	4590	),
(	4590	),
(	4590	),
(	4580	),
(	4580	),
(	4580	),
(	4580	),
(	4570	),
(	4570	),
(	4570	),
(	4560	),
(	4560	),
(	4560	),
(	4560	),
(	4550	),
(	4550	),
(	4550	),
(	4540	),
(	4540	),
(	4540	),
(	4530	),
(	4530	),
(	4530	),
(	4530	),
(	4520	),
(	4520	),
(	4520	),
(	4510	),
(	4510	),
(	4510	),
(	4510	),
(	4500	),
(	4500	),
(	4500	),
(	4490	),
(	4490	),
(	4490	),
(	4480	),
(	4480	),
(	4480	),
(	4480	),
(	4470	),
(	4470	),
(	4470	),
(	4460	),
(	4460	),
(	4460	),
(	4460	),
(	4450	),
(	4450	),
(	4450	),
(	4440	),
(	4440	),
(	4440	),
(	4430	),
(	4430	),
(	4430	),
(	4430	),
(	4420	),
(	4420	),
(	4420	),
(	4410	),
(	4410	),
(	4410	),
(	4410	),
(	4400	),
(	4400	),
(	4400	),
(	4390	),
(	4390	),
(	4390	),
(	4380	),
(	4380	),
(	4380	),
(	4380	),
(	4370	),
(	4370	),
(	4370	),
(	4360	),
(	4360	),
(	4360	),
(	4360	),
(	4350	),
(	4350	),
(	4350	),
(	4340	),
(	4340	),
(	4340	),
(	4330	),
(	4330	),
(	4330	),
(	4330	),
(	4320	),
(	4320	),
(	4320	),
(	4310	),
(	4310	),
(	4310	),
(	4310	),
(	4300	),
(	4300	),
(	4300	),
(	4290	),
(	4290	),
(	4290	),
(	4280	),
(	4280	),
(	4280	),
(	4280	),
(	4270	),
(	4270	),
(	4270	),
(	4260	),
(	4260	),
(	4260	),
(	4260	),
(	4250	),
(	4250	),
(	4250	),
(	4240	),
(	4240	),
(	4240	),
(	4230	),
(	4230	),
(	4230	),
(	4230	),
(	4220	),
(	4220	),
(	4220	),
(	4210	),
(	4210	),
(	4210	),
(	4210	),
(	4200	),
(	4200	),
(	4200	),
(	4190	),
(	4190	),
(	4190	),
(	4180	),
(	4180	),
(	4180	),
(	4180	),
(	4170	),
(	4170	),
(	4170	),
(	4160	),
(	4160	),
(	4160	),
(	4160	),
(	4150	),
(	4150	),
(	4150	),
(	4140	),
(	4140	),
(	4140	),
(	4130	),
(	4130	),
(	4130	),
(	4130	),
(	4120	),
(	4120	),
(	4120	),
(	4110	),
(	4110	),
(	4110	),
(	4110	),
(	4100	),
(	4100	),
(	4100	),
(	4090	),
(	4090	),
(	4090	),
(	4080	),
(	4080	),
(	4080	),
(	4080	),
(	4070	),
(	4070	),
(	4070	),
(	4060	),
(	4060	),
(	4060	),
(	4060	),
(	4050	),
(	4050	),
(	4050	),
(	4040	),
(	4040	),
(	4040	),
(	4030	),
(	4030	),
(	4030	),
(	4030	),
(	4020	),
(	4020	),
(	4020	),
(	4010	),
(	4010	),
(	4010	),
(	4010	),
(	4000	),
(	4000	),
(	4000	),
(	3990	),
(	3990	),
(	3990	),
(	3980	),
(	3980	),
(	3980	),
(	3980	),
(	3970	),
(	3970	),
(	3970	),
(	3960	),
(	3960	),
(	3960	),
(	3960	),
(	3950	),
(	3950	),
(	3950	),
(	3940	),
(	3940	),
(	3940	),
(	3930	),
(	3930	),
(	3930	),
(	3930	),
(	3920	),
(	3920	),
(	3920	),
(	3910	),
(	3910	),
(	3910	),
(	3910	),
(	3900	),
(	3900	),
(	3900	),
(	3890	),
(	3890	),
(	3890	),
(	3880	),
(	3880	),
(	3880	),
(	3880	),
(	3870	),
(	3870	),
(	3870	),
(	3860	),
(	3860	),
(	3860	),
(	3860	),
(	3850	),
(	3850	),
(	3850	),
(	3840	),
(	3840	),
(	3840	),
(	3830	),
(	3830	),
(	3830	),
(	3830	),
(	3820	),
(	3820	),
(	3820	),
(	3810	),
(	3810	),
(	3810	),
(	3810	),
(	3800	),
(	3800	),
(	3800	),
(	3790	),
(	3790	),
(	3790	),
(	3780	),
(	3780	),
(	3780	),
(	3780	),
(	3770	),
(	3770	),
(	3770	),
(	3760	),
(	3760	),
(	3760	),
(	3760	),
(	3750	),
(	3750	),
(	3750	),
(	3740	),
(	3740	),
(	3740	),
(	3730	),
(	3730	),
(	3730	),
(	3730	),
(	3720	),
(	3720	),
(	3720	),
(	3710	),
(	3710	),
(	3710	),
(	3710	),
(	3700	),
(	3700	),
(	3700	),
(	3690	),
(	3690	),
(	3690	),
(	3680	),
(	3680	),
(	3680	),
(	3680	),
(	3670	),
(	3670	),
(	3670	),
(	3660	),
(	3660	),
(	3660	),
(	3660	),
(	3650	),
(	3650	),
(	3650	),
(	3640	),
(	3640	),
(	3640	),
(	3630	),
(	3630	),
(	3630	),
(	3630	),
(	3620	),
(	3620	),
(	3620	),
(	3610	),
(	3610	),
(	3610	),
(	3610	),
(	3600	),
(	3600	),
(	3600	),
(	3590	),
(	3590	),
(	3590	),
(	3590	),
(	3580	),
(	3580	),
(	3580	),
(	3570	),
(	3570	),
(	3570	),
(	3560	),
(	3560	),
(	3560	),
(	3560	),
(	3550	),
(	3550	),
(	3550	),
(	3540	),
(	3540	),
(	3540	),
(	3540	),
(	3530	),
(	3530	),
(	3530	),
(	3520	),
(	3520	),
(	3520	),
(	3510	),
(	3510	),
(	3510	),
(	3510	),
(	3500	),
(	3500	),
(	3500	),
(	3490	),
(	3490	),
(	3490	),
(	3490	),
(	3480	),
(	3480	),
(	3480	),
(	3470	),
(	3470	),
(	3470	),
(	3460	),
(	3460	),
(	3460	),
(	3460	),
(	3450	),
(	3450	),
(	3450	),
(	3440	),
(	3440	),
(	3440	),
(	3440	),
(	3430	),
(	3430	),
(	3430	),
(	3420	),
(	3420	),
(	3420	),
(	3410	),
(	3410	),
(	3410	),
(	3410	),
(	3400	),
(	3400	),
(	3400	),
(	3390	),
(	3390	),
(	3390	),
(	3390	),
(	3380	),
(	3380	),
(	3380	),
(	3370	),
(	3370	),
(	3370	),
(	3360	),
(	3360	),
(	3360	),
(	3360	),
(	3350	),
(	3350	),
(	3350	),
(	3340	),
(	3340	),
(	3340	),
(	3340	),
(	3330	),
(	3330	),
(	3330	),
(	3320	),
(	3320	),
(	3320	),
(	3310	),
(	3310	),
(	3310	),
(	3310	),
(	3300	),
(	3300	),
(	3300	),
(	3290	),
(	3290	),
(	3290	),
(	3290	),
(	3280	),
(	3280	),
(	3280	),
(	3270	),
(	3270	),
(	3270	),
(	3260	),
(	3260	),
(	3260	),
(	3260	),
(	3250	),
(	3250	),
(	3250	),
(	3240	),
(	3240	),
(	3240	),
(	3240	),
(	3230	),
(	3230	),
(	3230	),
(	3220	),
(	3220	),
(	3220	),
(	3210	),
(	3210	),
(	3210	),
(	3210	),
(	3200	),
(	3200	),
(	3200	),
(	3190	),
(	3190	),
(	3190	),
(	3190	),
(	3180	),
(	3180	),
(	3180	),
(	3170	),
(	3170	),
(	3170	),
(	3160	),
(	3160	),
(	3160	),
(	3160	),
(	3150	),
(	3150	),
(	3150	),
(	3140	),
(	3140	),
(	3140	),
(	3140	),
(	3130	),
(	3130	),
(	3130	),
(	3120	),
(	3120	),
(	3120	),
(	3110	),
(	3110	),
(	3110	),
(	3110	),
(	3100	),
(	3100	),
(	3100	),
(	3090	),
(	3090	),
(	3090	),
(	3090	),
(	3080	),
(	3080	),
(	3080	),
(	3070	),
(	3070	),
(	3070	),
(	3060	),
(	3060	),
(	3060	),
(	3060	),
(	3050	),
(	3050	),
(	3050	),
(	3040	),
(	3040	),
(	3040	),
(	3040	),
(	3030	),
(	3030	),
(	3030	),
(	3020	),
(	3020	),
(	3020	),
(	3010	),
(	3010	),
(	3010	),
(	3010	),
(	3000	),
(	3000	),
(	3000	),
(	2990	),
(	2990	),
(	2990	),
(	2990	),
(	2980	),
(	2980	),
(	2980	),
(	2970	),
(	2970	),
(	2970	),
(	2960	),
(	2960	),
(	2960	),
(	2960	),
(	2950	),
(	2950	),
(	2950	),
(	2940	),
(	2940	),
(	2940	),
(	2940	),
(	2930	),
(	2930	),
(	2930	),
(	2920	),
(	2920	),
(	2920	),
(	2910	),
(	2910	),
(	2910	),
(	2910	),
(	2900	),
(	2900	),
(	2900	),
(	2890	),
(	2890	),
(	2890	),
(	2890	),
(	2880	),
(	2880	),
(	2880	),
(	2870	),
(	2870	),
(	2870	),
(	2860	),
(	2860	),
(	2860	),
(	2860	),
(	2850	),
(	2850	),
(	2850	),
(	2840	),
(	2840	),
(	2840	),
(	2840	),
(	2830	),
(	2830	),
(	2830	),
(	2820	),
(	2820	),
(	2820	),
(	2810	),
(	2810	),
(	2810	),
(	2810	),
(	2800	),
(	2800	),
(	2800	),
(	2790	),
(	2790	),
(	2790	),
(	2790	),
(	2780	),
(	2780	),
(	2780	),
(	2770	),
(	2770	),
(	2770	),
(	2760	),
(	2760	),
(	2760	),
(	2760	),
(	2750	),
(	2750	),
(	2750	),
(	2740	),
(	2740	),
(	2740	),
(	2740	),
(	2730	),
(	2730	),
(	2730	),
(	2720	),
(	2720	),
(	2720	),
(	2710	),
(	2710	),
(	2710	),
(	2710	),
(	2700	),
(	2700	),
(	2700	),
(	2690	),
(	2690	),
(	2690	),
(	2690	),
(	2680	),
(	2680	),
(	2680	),
(	2670	),
(	2670	),
(	2670	),
(	2660	),
(	2660	),
(	2660	),
(	2660	),
(	2650	),
(	2650	),
(	2650	),
(	2640	),
(	2640	),
(	2640	),
(	2640	),
(	2630	),
(	2630	),
(	2630	),
(	2620	),
(	2620	),
(	2620	),
(	2610	),
(	2610	),
(	2610	),
(	2610	),
(	2600	),
(	2600	),
(	2600	),
(	2590	),
(	2590	),
(	2590	),
(	2590	),
(	2580	),
(	2580	),
(	2580	),
(	2570	),
(	2570	),
(	2570	),
(	2560	),
(	2560	),
(	2560	),
(	2560	),
(	2550	),
(	2550	),
(	2550	),
(	2540	),
(	2540	),
(	2540	),
(	2540	),
(	2530	),
(	2530	),
(	2530	),
(	2520	),
(	2520	),
(	2520	),
(	2510	),
(	2510	),
(	2510	),
(	2510	),
(	2500	),
(	2500	),
(	2500	),
(	2490	),
(	2490	),
(	2490	),
(	2490	),
(	2480	),
(	2480	),
(	2480	),
(	2470	),
(	2470	),
(	2470	),
(	2460	),
(	2460	),
(	2460	),
(	2460	),
(	2450	),
(	2450	),
(	2450	),
(	2440	),
(	2440	),
(	2440	),
(	2440	),
(	2430	),
(	2430	),
(	2430	),
(	2420	),
(	2420	),
(	2420	),
(	2410	),
(	2410	),
(	2410	),
(	2410	),
(	2400	),
(	2400	),
(	2400	),
(	2390	),
(	2390	),
(	2390	),
(	2390	),
(	2380	),
(	2380	),
(	2380	),
(	2370	),
(	2370	),
(	2370	),
(	2360	),
(	2360	),
(	2360	),
(	2360	),
(	2350	),
(	2350	),
(	2350	),
(	2340	),
(	2340	),
(	2340	),
(	2340	),
(	2330	),
(	2330	),
(	2330	),
(	2320	),
(	2320	),
(	2320	),
(	2310	),
(	2310	),
(	2310	),
(	2310	),
(	2300	),
(	2300	),
(	2300	),
(	2290	),
(	2290	),
(	2290	),
(	2290	),
(	2280	),
(	2280	),
(	2280	),
(	2270	),
(	2270	),
(	2270	),
(	2260	),
(	2260	),
(	2260	),
(	2260	),
(	2250	),
(	2250	),
(	2250	),
(	2240	),
(	2240	),
(	2240	),
(	2240	),
(	2230	),
(	2230	),
(	2230	),
(	2220	),
(	2220	),
(	2220	),
(	2220	),
(	2210	),
(	2210	),
(	2210	),
(	2200	),
(	2200	),
(	2200	),
(	2190	),
(	2190	),
(	2190	),
(	2190	),
(	2180	),
(	2180	),
(	2180	),
(	2170	),
(	2170	),
(	2170	),
(	2170	),
(	2160	),
(	2160	),
(	2160	),
(	2150	),
(	2150	),
(	2150	),
(	2140	),
(	2140	),
(	2140	),
(	2140	),
(	2130	),
(	2130	),
(	2130	),
(	2120	),
(	2120	),
(	2120	),
(	2120	),
(	2110	),
(	2110	),
(	2110	),
(	2100	),
(	2100	),
(	2100	),
(	2090	),
(	2090	),
(	2090	),
(	2090	),
(	2080	),
(	2080	),
(	2080	),
(	2070	),
(	2070	),
(	2070	),
(	2070	),
(	2060	),
(	2060	),
(	2060	),
(	2050	),
(	2050	),
(	2050	),
(	2040	),
(	2040	),
(	2040	),
(	2040	),
(	2030	),
(	2030	),
(	2030	),
(	2020	),
(	2020	),
(	2020	),
(	2020	),
(	2010	),
(	2010	),
(	2010	),
(	2000	),
(	2000	),
(	2000	),
(	1990	),
(	1990	),
(	1990	),
(	1990	),
(	1980	),
(	1980	),
(	1980	),
(	1970	),
(	1970	),
(	1970	),
(	1970	),
(	1960	),
(	1960	),
(	1960	),
(	1950	),
(	1950	),
(	1950	),
(	1940	),
(	1940	),
(	1940	),
(	1940	),
(	1930	),
(	1930	),
(	1930	),
(	1920	),
(	1920	),
(	1920	),
(	1920	),
(	1910	),
(	1910	),
(	1910	),
(	1900	),
(	1900	),
(	1900	),
(	1890	),
(	1890	),
(	1890	),
(	1890	),
(	1880	),
(	1880	),
(	1880	),
(	1870	),
(	1870	),
(	1870	),
(	1870	),
(	1860	),
(	1860	),
(	1860	),
(	1850	),
(	1850	),
(	1850	),
(	1840	),
(	1840	),
(	1840	),
(	1840	),
(	1830	),
(	1830	),
(	1830	),
(	1820	),
(	1820	),
(	1820	),
(	1820	),
(	1810	),
(	1810	),
(	1810	),
(	1800	),
(	1800	),
(	1800	),
(	1790	),
(	1790	),
(	1790	),
(	1790	),
(	1780	),
(	1780	),
(	1780	),
(	1770	),
(	1770	),
(	1770	),
(	1770	),
(	1760	),
(	1760	),
(	1760	),
(	1750	),
(	1750	),
(	1750	),
(	1740	),
(	1740	),
(	1740	),
(	1740	),
(	1730	),
(	1730	),
(	1730	),
(	1720	),
(	1720	),
(	1720	),
(	1720	),
(	1710	),
(	1710	),
(	1710	),
(	1700	),
(	1700	),
(	1700	),
(	1690	),
(	1690	),
(	1690	),
(	1690	),
(	1680	),
(	1680	),
(	1680	),
(	1670	),
(	1670	),
(	1670	),
(	1670	),
(	1660	),
(	1660	),
(	1660	),
(	1650	),
(	1650	),
(	1650	),
(	1640	),
(	1640	),
(	1640	),
(	1640	),
(	1630	),
(	1630	),
(	1630	),
(	1620	),
(	1620	),
(	1620	),
(	1620	),
(	1610	),
(	1610	),
(	1610	),
(	1600	),
(	1600	),
(	1600	),
(	1590	),
(	1590	),
(	1590	),
(	1590	),
(	1580	),
(	1580	),
(	1580	),
(	1570	),
(	1570	),
(	1570	),
(	1570	),
(	1560	),
(	1560	),
(	1560	),
(	1550	),
(	1550	),
(	1550	),
(	1540	),
(	1540	),
(	1540	),
(	1540	),
(	1530	),
(	1530	),
(	1530	),
(	1520	),
(	1520	),
(	1520	),
(	1520	),
(	1510	),
(	1510	),
(	1510	),
(	1500	),
(	1500	),
(	1500	),
(	1490	),
(	1490	),
(	1490	),
(	1490	),
(	1480	),
(	1480	),
(	1480	),
(	1470	),
(	1470	),
(	1470	),
(	1470	),
(	1460	),
(	1460	),
(	1460	),
(	1450	),
(	1450	),
(	1450	),
(	1440	),
(	1440	),
(	1440	),
(	1440	),
(	1430	),
(	1430	),
(	1430	),
(	1420	),
(	1420	),
(	1420	),
(	1420	),
(	1410	),
(	1410	),
(	1410	),
(	1400	),
(	1400	),
(	1400	),
(	1390	),
(	1390	),
(	1390	),
(	1390	),
(	1380	),
(	1380	),
(	1380	),
(	1370	),
(	1370	),
(	1370	),
(	1370	),
(	1360	),
(	1360	),
(	1360	),
(	1350	),
(	1350	),
(	1350	),
(	1340	),
(	1340	),
(	1340	),
(	1340	),
(	1330	),
(	1330	),
(	1330	),
(	1320	),
(	1320	),
(	1320	),
(	1320	),
(	1310	),
(	1310	),
(	1310	),
(	1300	),
(	1300	),
(	1300	),
(	1290	),
(	1290	),
(	1290	),
(	1290	),
(	1280	),
(	1280	),
(	1280	),
(	1270	),
(	1270	),
(	1270	),
(	1270	),
(	1260	),
(	1260	),
(	1260	),
(	1250	),
(	1250	),
(	1250	),
(	1240	),
(	1240	),
(	1240	),
(	1240	),
(	1230	),
(	1230	),
(	1230	),
(	1220	),
(	1220	),
(	1220	),
(	1220	),
(	1210	),
(	1210	),
(	1210	),
(	1200	),
(	1200	),
(	1200	),
(	1190	),
(	1190	),
(	1190	),
(	1190	),
(	1180	),
(	1180	),
(	1180	),
(	1170	),
(	1170	),
(	1170	),
(	1170	),
(	1160	),
(	1160	),
(	1160	),
(	1150	),
(	1150	),
(	1150	),
(	1140	),
(	1140	),
(	1140	),
(	1140	),
(	1130	),
(	1130	),
(	1130	),
(	1120	),
(	1120	),
(	1120	),
(	1120	),
(	1110	),
(	1110	),
(	1110	),
(	1100	),
(	1100	),
(	1100	),
(	1090	),
(	1090	),
(	1090	),
(	1090	),
(	1080	),
(	1080	),
(	1080	),
(	1070	),
(	1070	),
(	1070	),
(	1070	),
(	1060	),
(	1060	),
(	1060	),
(	1050	),
(	1050	),
(	1050	),
(	1040	),
(	1040	),
(	1040	),
(	1040	),
(	1030	),
(	1030	),
(	1030	),
(	1020	),
(	1020	),
(	1020	),
(	1020	),
(	1010	),
(	1010	),
(	1010	),
(	1000	),
(	1000	),
(	1000	),
(	990	),
(	990	),
(	990	),
(	990	),
(	980	),
(	980	),
(	980	),
(	970	),
(	970	),
(	970	),
(	970	),
(	960	),
(	960	),
(	960	),
(	950	),
(	950	),
(	950	),
(	940	),
(	940	),
(	940	),
(	940	),
(	930	),
(	930	),
(	930	),
(	920	),
(	920	),
(	920	),
(	920	),
(	910	),
(	910	),
(	910	),
(	900	),
(	900	),
(	900	),
(	890	),
(	890	),
(	890	),
(	890	),
(	880	),
(	880	),
(	880	),
(	870	),
(	870	),
(	870	),
(	870	),
(	860	),
(	860	),
(	860	),
(	850	),
(	850	),
(	850	),
(	850	),
(	840	),
(	840	),
(	840	),
(	830	),
(	830	),
(	830	),
(	820	),
(	820	),
(	820	),
(	820	),
(	810	),
(	810	),
(	810	),
(	800	),
(	800	),
(	800	),
(	800	),
(	790	),
(	790	),
(	790	),
(	780	),
(	780	),
(	780	),
(	770	),
(	770	),
(	770	),
(	770	),
(	760	),
(	760	),
(	760	),
(	750	),
(	750	),
(	750	),
(	750	),
(	740	),
(	740	),
(	740	),
(	730	),
(	730	),
(	730	),
(	720	),
(	720	),
(	720	),
(	720	),
(	710	),
(	710	),
(	710	),
(	700	),
(	700	),
(	700	),
(	700	),
(	690	),
(	690	),
(	690	),
(	680	),
(	680	),
(	680	),
(	670	),
(	670	),
(	670	),
(	670	),
(	660	),
(	660	),
(	660	),
(	650	),
(	650	),
(	650	),
(	650	),
(	640	),
(	640	),
(	640	),
(	630	),
(	630	),
(	630	),
(	620	),
(	620	),
(	620	),
(	620	),
(	610	),
(	610	),
(	610	),
(	600	),
(	600	),
(	600	),
(	600	),
(	590	),
(	590	),
(	590	),
(	580	),
(	580	),
(	580	),
(	570	),
(	570	),
(	570	),
(	570	),
(	560	),
(	560	),
(	560	),
(	550	),
(	550	),
(	550	),
(	550	),
(	540	),
(	540	),
(	540	),
(	530	),
(	530	),
(	530	),
(	520	),
(	520	),
(	520	),
(	520	),
(	510	),
(	510	),
(	510	),
(	500	),
(	500	),
(	500	),
(	500	),
(	490	),
(	490	),
(	490	),
(	480	),
(	480	),
(	480	),
(	470	),
(	470	),
(	470	),
(	470	),
(	460	),
(	460	),
(	460	),
(	450	),
(	450	),
(	450	),
(	450	),
(	440	),
(	440	),
(	440	),
(	430	),
(	430	),
(	430	),
(	420	),
(	420	),
(	420	),
(	420	),
(	410	),
(	410	),
(	410	),
(	400	),
(	400	),
(	400	),
(	400	),
(	390	),
(	390	),
(	390	),
(	380	),
(	380	),
(	380	),
(	370	),
(	370	),
(	370	),
(	370	),
(	360	),
(	360	),
(	360	),
(	350	),
(	350	),
(	350	),
(	350	),
(	340	),
(	340	),
(	340	),
(	330	),
(	330	),
(	330	),
(	320	),
(	320	),
(	320	),
(	320	),
(	310	),
(	310	),
(	310	),
(	300	),
(	300	),
(	300	),
(	300	),
(	290	),
(	290	),
(	290	),
(	280	),
(	280	),
(	280	),
(	270	),
(	270	),
(	270	),
(	270	),
(	260	),
(	260	),
(	260	),
(	250	),
(	250	),
(	250	),
(	250	),
(	240	),
(	240	),
(	240	),
(	230	),
(	230	),
(	230	),
(	220	),
(	220	),
(	220	),
(	220	),
(	210	),
(	210	),
(	210	),
(	200	),
(	200	),
(	200	),
(	200	),
(	190	),
(	190	),
(	190	),
(	180	),
(	180	),
(	180	),
(	170	),
(	170	),
(	170	),
(	170	),
(	160	),
(	160	),
(	160	),
(	150	),
(	150	),
(	150	),
(	150	),
(	140	),
(	140	),
(	140	),
(	130	),
(	130	),
(	130	),
(	120	),
(	120	),
(	120	),
(	120	),
(	110	),
(	110	),
(	110	),
(	100	),
(	100	),
(	100	),
(	100	),
(	90	),
(	90	),
(	90	),
(	80	),
(	80	),
(	80	),
(	70	),
(	70	),
(	70	),
(	70	),
(	60	),
(	60	),
(	60	),
(	50	),
(	50	),
(	50	),
(	50	),
(	40	),
(	40	),
(	40	),
(	30	),
(	30	),
(	30	),
(	20	),
(	20	),
(	20	),
(	20	),
(	10	),
(	10	),
(	10	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	),
(	0	)
);
begin

cycle <= std_logic_vector(to_unsigned(d2c_LUT(to_integer(unsigned(distance))),cycle'length));
							
end behavior;